package rbr_pkg;

typedef struct packed{
    logic   plus;
    logic   minus;
}  signed_digit;


endpackage